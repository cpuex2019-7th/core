y0n3uchy@y0n3uchy.local.1211