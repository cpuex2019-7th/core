`default_nettype none

module uart_buffer(
	               input wire         clk,
	               input wire         rstn,

	               // Bus for MMU
                   ////////////
	               input wire [3:0]   mmu_axi_araddr,
	               output reg         mmu_axi_arready,
	               input wire         mmu_axi_arvalid,
	               input wire [2:0]   mmu_axi_arprot, 

	               input wire         mmu_axi_bready,
	               output wire [1:0]  mmu_axi_bresp,
	               output wire        mmu_axi_bvalid,

	               output reg [31:0]  mmu_axi_rdata,
	               input wire         mmu_axi_rready,
	               output reg [1:0]   mmu_axi_rresp,
	               output reg         mmu_axi_rvalid,

	               input wire [3:0]   mmu_axi_awaddr,
	               output wire        mmu_axi_awready,
	               input wire         mmu_axi_awvalid,
	               input wire [2:0]   mmu_axi_awprot, 

	               input wire [31:0]  mmu_axi_wdata,
	               output wire        mmu_axi_wready,
	               input wire [3:0]   mmu_axi_wstrb,
	               input wire         mmu_axi_wvalid,

                   // Bus for UART
                   ////////////
	               output reg [3:0]   uart_axi_araddr,
	               input wire         uart_axi_arready,
	               output reg         uart_axi_arvalid,
	               output reg [2:0]   uart_axi_arprot, 

                   // response channel
	               output wire        uart_axi_bready,
	               input wire [1:0]   uart_axi_bresp,
	               input wire         uart_axi_bvalid,

                   // read data channel
	               input wire [31:0]  uart_axi_rdata,
	               output reg         uart_axi_rready,
	               input wire [1:0]   uart_axi_rresp,
	               input wire         uart_axi_rvalid,

                   // address write channel
	               output wire [3:0]  uart_axi_awaddr,
	               input wire         uart_axi_awready,
	               output wire        uart_axi_awvalid,
	               output wire [2:0]  uart_axi_awprot, 

                   // data write channel
	               output wire [31:0] uart_axi_wdata,
	               input wire         uart_axi_wready,
	               output wire [3:0]  uart_axi_wstrb,
	               output wire        uart_axi_wvalid);

   // bypass wires related to uart tx
   assign mmu_axi_bready = uart_axi_bready;
   assign uart_axi_bresp = mmu_axi_bresp;
   assign uart_axi_bvalid = mmu_axi_bvalid;
   
   assign uart_axi_awaddr = mmu_axi_awaddr;
   assign mmu_axi_awready = uart_axi_awready;
   assign  uart_axi_awvalid = mmu_axi_awvalid;
   assign uart_axi_awprot = mmu_axi_awprot;

   assign uart_axi_wdata = mmu_axi_wdata;
   assign mmu_axi_wready = uart_axi_wready;
   assign uart_axi_wstrb = mmu_axi_wstrb;
   assign uart_axi_wvalid = mmu_axi_wvalid;
   

   reg [3:0]                          reading_state;
   localparam r_waiting_ready = 0;   
   localparam r_writing_ready = 1;   
   localparam r_waiting_data = 2;   
   localparam r_writing_data = 3;
   localparam r_waiting_uartlite_arready = 4;
   localparam r_waiting_uartlite_rvalid = 5;
   
   
   reg [7:0]                          buffer[2048];
   (* mark_debug = "true" *) reg [10:0]   head_idx;
   (* mark_debug = "true" *) reg [10:0]   tail_idx;
   (* mark_debug = "true" *)  wire         is_buffer_empty = (tail_idx - head_idx == 0);
   
   initial begin
      mmu_axi_arready <= 1;
      mmu_axi_rvalid <= 0;
      
      uart_axi_arvalid <= 0;
      uart_axi_rready <= 0;

      head_idx <= 0;
      tail_idx <= 1300;
      
      reading_state <= r_waiting_ready;      

      buffer[0] = 8'd194;
      buffer[1] = 8'd140;
      buffer[2] = 8'd0;
      buffer[3] = 8'd0;
      buffer[4] = 8'd66;
      buffer[5] = 8'd12;
      buffer[6] = 8'd0;
      buffer[7] = 8'd0;
      buffer[8] = 8'd193;
      buffer[9] = 8'd160;
      buffer[10] = 8'd0;
      buffer[11] = 8'd0;
      buffer[12] = 8'd65;
      buffer[13] = 8'd160;
      buffer[14] = 8'd0;
      buffer[15] = 8'd0;
      buffer[16] = 8'd65;
      buffer[17] = 8'd240;
      buffer[18] = 8'd0;
      buffer[19] = 8'd0;
      buffer[20] = 8'd63;
      buffer[21] = 8'd128;
      buffer[22] = 8'd0;
      buffer[23] = 8'd0;
      buffer[24] = 8'd66;
      buffer[25] = 8'd72;
      buffer[26] = 8'd0;
      buffer[27] = 8'd0;
      buffer[28] = 8'd66;
      buffer[29] = 8'd72;
      buffer[30] = 8'd0;
      buffer[31] = 8'd0;
      buffer[32] = 8'd67;
      buffer[33] = 8'd127;
      buffer[34] = 8'd0;
      buffer[35] = 8'd0;
      buffer[36] = 8'd0;
      buffer[37] = 8'd0;
      buffer[38] = 8'd0;
      buffer[39] = 8'd0;
      buffer[40] = 8'd0;
      buffer[41] = 8'd0;
      buffer[42] = 8'd0;
      buffer[43] = 8'd1;
      buffer[44] = 8'd0;
      buffer[45] = 8'd0;
      buffer[46] = 8'd0;
      buffer[47] = 8'd1;
      buffer[48] = 8'd0;
      buffer[49] = 8'd0;
      buffer[50] = 8'd0;
      buffer[51] = 8'd0;
      buffer[52] = 8'd65;
      buffer[53] = 8'd160;
      buffer[54] = 8'd0;
      buffer[55] = 8'd0;
      buffer[56] = 8'd65;
      buffer[57] = 8'd160;
      buffer[58] = 8'd0;
      buffer[59] = 8'd0;
      buffer[60] = 8'd66;
      buffer[61] = 8'd130;
      buffer[62] = 8'd0;
      buffer[63] = 8'd0;
      buffer[64] = 8'd0;
      buffer[65] = 8'd0;
      buffer[66] = 8'd0;
      buffer[67] = 8'd0;
      buffer[68] = 8'd65;
      buffer[69] = 8'd160;
      buffer[70] = 8'd0;
      buffer[71] = 8'd0;
      buffer[72] = 8'd66;
      buffer[73] = 8'd52;
      buffer[74] = 8'd0;
      buffer[75] = 8'd0;
      buffer[76] = 8'd63;
      buffer[77] = 8'd128;
      buffer[78] = 8'd0;
      buffer[79] = 8'd0;
      buffer[80] = 8'd63;
      buffer[81] = 8'd128;
      buffer[82] = 8'd0;
      buffer[83] = 8'd0;
      buffer[84] = 8'd67;
      buffer[85] = 8'd122;
      buffer[86] = 8'd0;
      buffer[87] = 8'd0;
      buffer[88] = 8'd67;
      buffer[89] = 8'd0;
      buffer[90] = 8'd0;
      buffer[91] = 8'd0;
      buffer[92] = 8'd67;
      buffer[93] = 8'd82;
      buffer[94] = 8'd0;
      buffer[95] = 8'd0;
      buffer[96] = 8'd0;
      buffer[97] = 8'd0;
      buffer[98] = 8'd0;
      buffer[99] = 8'd0;
      buffer[100] = 8'd0;
      buffer[101] = 8'd0;
      buffer[102] = 8'd0;
      buffer[103] = 8'd0;
      buffer[104] = 8'd0;
      buffer[105] = 8'd0;
      buffer[106] = 8'd0;
      buffer[107] = 8'd3;
      buffer[108] = 8'd0;
      buffer[109] = 8'd0;
      buffer[110] = 8'd0;
      buffer[111] = 8'd1;
      buffer[112] = 8'd0;
      buffer[113] = 8'd0;
      buffer[114] = 8'd0;
      buffer[115] = 8'd0;
      buffer[116] = 8'd65;
      buffer[117] = 8'd200;
      buffer[118] = 8'd0;
      buffer[119] = 8'd0;
      buffer[120] = 8'd66;
      buffer[121] = 8'd32;
      buffer[122] = 8'd0;
      buffer[123] = 8'd0;
      buffer[124] = 8'd66;
      buffer[125] = 8'd140;
      buffer[126] = 8'd0;
      buffer[127] = 8'd0;
      buffer[128] = 8'd0;
      buffer[129] = 8'd0;
      buffer[130] = 8'd0;
      buffer[131] = 8'd0;
      buffer[132] = 8'd0;
      buffer[133] = 8'd0;
      buffer[134] = 8'd0;
      buffer[135] = 8'd0;
      buffer[136] = 8'd66;
      buffer[137] = 8'd32;
      buffer[138] = 8'd0;
      buffer[139] = 8'd0;
      buffer[140] = 8'd63;
      buffer[141] = 8'd128;
      buffer[142] = 8'd0;
      buffer[143] = 8'd0;
      buffer[144] = 8'd63;
      buffer[145] = 8'd128;
      buffer[146] = 8'd0;
      buffer[147] = 8'd0;
      buffer[148] = 8'd67;
      buffer[149] = 8'd122;
      buffer[150] = 8'd0;
      buffer[151] = 8'd0;
      buffer[152] = 8'd67;
      buffer[153] = 8'd0;
      buffer[154] = 8'd0;
      buffer[155] = 8'd0;
      buffer[156] = 8'd67;
      buffer[157] = 8'd82;
      buffer[158] = 8'd0;
      buffer[159] = 8'd0;
      buffer[160] = 8'd0;
      buffer[161] = 8'd0;
      buffer[162] = 8'd0;
      buffer[163] = 8'd0;
      buffer[164] = 8'd0;
      buffer[165] = 8'd0;
      buffer[166] = 8'd0;
      buffer[167] = 8'd0;
      buffer[168] = 8'd0;
      buffer[169] = 8'd0;
      buffer[170] = 8'd0;
      buffer[171] = 8'd3;
      buffer[172] = 8'd0;
      buffer[173] = 8'd0;
      buffer[174] = 8'd0;
      buffer[175] = 8'd1;
      buffer[176] = 8'd0;
      buffer[177] = 8'd0;
      buffer[178] = 8'd0;
      buffer[179] = 8'd0;
      buffer[180] = 8'd0;
      buffer[181] = 8'd0;
      buffer[182] = 8'd0;
      buffer[183] = 8'd0;
      buffer[184] = 8'd65;
      buffer[185] = 8'd240;
      buffer[186] = 8'd0;
      buffer[187] = 8'd0;
      buffer[188] = 8'd65;
      buffer[189] = 8'd240;
      buffer[190] = 8'd0;
      buffer[191] = 8'd0;
      buffer[192] = 8'd0;
      buffer[193] = 8'd0;
      buffer[194] = 8'd0;
      buffer[195] = 8'd0;
      buffer[196] = 8'd192;
      buffer[197] = 8'd160;
      buffer[198] = 8'd0;
      buffer[199] = 8'd0;
      buffer[200] = 8'd0;
      buffer[201] = 8'd0;
      buffer[202] = 8'd0;
      buffer[203] = 8'd0;
      buffer[204] = 8'd191;
      buffer[205] = 8'd128;
      buffer[206] = 8'd0;
      buffer[207] = 8'd0;
      buffer[208] = 8'd63;
      buffer[209] = 8'd128;
      buffer[210] = 8'd0;
      buffer[211] = 8'd0;
      buffer[212] = 8'd67;
      buffer[213] = 8'd122;
      buffer[214] = 8'd0;
      buffer[215] = 8'd0;
      buffer[216] = 8'd67;
      buffer[217] = 8'd0;
      buffer[218] = 8'd0;
      buffer[219] = 8'd0;
      buffer[220] = 8'd67;
      buffer[221] = 8'd83;
      buffer[222] = 8'd0;
      buffer[223] = 8'd0;
      buffer[224] = 8'd0;
      buffer[225] = 8'd0;
      buffer[226] = 8'd0;
      buffer[227] = 8'd0;
      buffer[228] = 8'd0;
      buffer[229] = 8'd0;
      buffer[230] = 8'd0;
      buffer[231] = 8'd0;
      buffer[232] = 8'd0;
      buffer[233] = 8'd0;
      buffer[234] = 8'd0;
      buffer[235] = 8'd1;
      buffer[236] = 8'd0;
      buffer[237] = 8'd0;
      buffer[238] = 8'd0;
      buffer[239] = 8'd1;
      buffer[240] = 8'd0;
      buffer[241] = 8'd0;
      buffer[242] = 8'd0;
      buffer[243] = 8'd0;
      buffer[244] = 8'd65;
      buffer[245] = 8'd160;
      buffer[246] = 8'd0;
      buffer[247] = 8'd0;
      buffer[248] = 8'd65;
      buffer[249] = 8'd32;
      buffer[250] = 8'd0;
      buffer[251] = 8'd0;
      buffer[252] = 8'd65;
      buffer[253] = 8'd240;
      buffer[254] = 8'd0;
      buffer[255] = 8'd0;
      buffer[256] = 8'd0;
      buffer[257] = 8'd0;
      buffer[258] = 8'd0;
      buffer[259] = 8'd0;
      buffer[260] = 8'd193;
      buffer[261] = 8'd32;
      buffer[262] = 8'd0;
      buffer[263] = 8'd0;
      buffer[264] = 8'd66;
      buffer[265] = 8'd160;
      buffer[266] = 8'd0;
      buffer[267] = 8'd0;
      buffer[268] = 8'd63;
      buffer[269] = 8'd128;
      buffer[270] = 8'd0;
      buffer[271] = 8'd0;
      buffer[272] = 8'd63;
      buffer[273] = 8'd128;
      buffer[274] = 8'd0;
      buffer[275] = 8'd0;
      buffer[276] = 8'd67;
      buffer[277] = 8'd122;
      buffer[278] = 8'd0;
      buffer[279] = 8'd0;
      buffer[280] = 8'd67;
      buffer[281] = 8'd0;
      buffer[282] = 8'd0;
      buffer[283] = 8'd0;
      buffer[284] = 8'd67;
      buffer[285] = 8'd83;
      buffer[286] = 8'd0;
      buffer[287] = 8'd0;
      buffer[288] = 8'd0;
      buffer[289] = 8'd0;
      buffer[290] = 8'd0;
      buffer[291] = 8'd0;
      buffer[292] = 8'd0;
      buffer[293] = 8'd0;
      buffer[294] = 8'd0;
      buffer[295] = 8'd0;
      buffer[296] = 8'd0;
      buffer[297] = 8'd0;
      buffer[298] = 8'd0;
      buffer[299] = 8'd2;
      buffer[300] = 8'd0;
      buffer[301] = 8'd0;
      buffer[302] = 8'd0;
      buffer[303] = 8'd1;
      buffer[304] = 8'd0;
      buffer[305] = 8'd0;
      buffer[306] = 8'd0;
      buffer[307] = 8'd0;
      buffer[308] = 8'd0;
      buffer[309] = 8'd0;
      buffer[310] = 8'd0;
      buffer[311] = 8'd0;
      buffer[312] = 8'd191;
      buffer[313] = 8'd192;
      buffer[314] = 8'd0;
      buffer[315] = 8'd0;
      buffer[316] = 8'd191;
      buffer[317] = 8'd128;
      buffer[318] = 8'd0;
      buffer[319] = 8'd0;
      buffer[320] = 8'd0;
      buffer[321] = 8'd0;
      buffer[322] = 8'd0;
      buffer[323] = 8'd0;
      buffer[324] = 8'd0;
      buffer[325] = 8'd0;
      buffer[326] = 8'd0;
      buffer[327] = 8'd0;
      buffer[328] = 8'd66;
      buffer[329] = 8'd72;
      buffer[330] = 8'd0;
      buffer[331] = 8'd0;
      buffer[332] = 8'd63;
      buffer[333] = 8'd128;
      buffer[334] = 8'd0;
      buffer[335] = 8'd0;
      buffer[336] = 8'd63;
      buffer[337] = 8'd128;
      buffer[338] = 8'd0;
      buffer[339] = 8'd0;
      buffer[340] = 8'd67;
      buffer[341] = 8'd122;
      buffer[342] = 8'd0;
      buffer[343] = 8'd0;
      buffer[344] = 8'd67;
      buffer[345] = 8'd0;
      buffer[346] = 8'd0;
      buffer[347] = 8'd0;
      buffer[348] = 8'd67;
      buffer[349] = 8'd83;
      buffer[350] = 8'd0;
      buffer[351] = 8'd0;
      buffer[352] = 8'd0;
      buffer[353] = 8'd0;
      buffer[354] = 8'd0;
      buffer[355] = 8'd0;
      buffer[356] = 8'd0;
      buffer[357] = 8'd0;
      buffer[358] = 8'd0;
      buffer[359] = 8'd0;
      buffer[360] = 8'd0;
      buffer[361] = 8'd0;
      buffer[362] = 8'd0;
      buffer[363] = 8'd1;
      buffer[364] = 8'd0;
      buffer[365] = 8'd0;
      buffer[366] = 8'd0;
      buffer[367] = 8'd1;
      buffer[368] = 8'd0;
      buffer[369] = 8'd0;
      buffer[370] = 8'd0;
      buffer[371] = 8'd0;
      buffer[372] = 8'd65;
      buffer[373] = 8'd176;
      buffer[374] = 8'd0;
      buffer[375] = 8'd0;
      buffer[376] = 8'd65;
      buffer[377] = 8'd224;
      buffer[378] = 8'd0;
      buffer[379] = 8'd0;
      buffer[380] = 8'd65;
      buffer[381] = 8'd224;
      buffer[382] = 8'd0;
      buffer[383] = 8'd0;
      buffer[384] = 8'd0;
      buffer[385] = 8'd0;
      buffer[386] = 8'd0;
      buffer[387] = 8'd0;
      buffer[388] = 8'd192;
      buffer[389] = 8'd160;
      buffer[390] = 8'd0;
      buffer[391] = 8'd0;
      buffer[392] = 8'd0;
      buffer[393] = 8'd0;
      buffer[394] = 8'd0;
      buffer[395] = 8'd0;
      buffer[396] = 8'd63;
      buffer[397] = 8'd128;
      buffer[398] = 8'd0;
      buffer[399] = 8'd0;
      buffer[400] = 8'd63;
      buffer[401] = 8'd128;
      buffer[402] = 8'd0;
      buffer[403] = 8'd0;
      buffer[404] = 8'd67;
      buffer[405] = 8'd122;
      buffer[406] = 8'd0;
      buffer[407] = 8'd0;
      buffer[408] = 8'd0;
      buffer[409] = 8'd0;
      buffer[410] = 8'd0;
      buffer[411] = 8'd0;
      buffer[412] = 8'd67;
      buffer[413] = 8'd83;
      buffer[414] = 8'd0;
      buffer[415] = 8'd0;
      buffer[416] = 8'd67;
      buffer[417] = 8'd83;
      buffer[418] = 8'd0;
      buffer[419] = 8'd0;
      buffer[420] = 8'd0;
      buffer[421] = 8'd0;
      buffer[422] = 8'd0;
      buffer[423] = 8'd0;
      buffer[424] = 8'd0;
      buffer[425] = 8'd0;
      buffer[426] = 8'd0;
      buffer[427] = 8'd3;
      buffer[428] = 8'd0;
      buffer[429] = 8'd0;
      buffer[430] = 8'd0;
      buffer[431] = 8'd1;
      buffer[432] = 8'd0;
      buffer[433] = 8'd0;
      buffer[434] = 8'd0;
      buffer[435] = 8'd0;
      buffer[436] = 8'd66;
      buffer[437] = 8'd32;
      buffer[438] = 8'd0;
      buffer[439] = 8'd0;
      buffer[440] = 8'd65;
      buffer[441] = 8'd224;
      buffer[442] = 8'd0;
      buffer[443] = 8'd0;
      buffer[444] = 8'd65;
      buffer[445] = 8'd224;
      buffer[446] = 8'd0;
      buffer[447] = 8'd0;
      buffer[448] = 8'd0;
      buffer[449] = 8'd0;
      buffer[450] = 8'd0;
      buffer[451] = 8'd0;
      buffer[452] = 8'd192;
      buffer[453] = 8'd160;
      buffer[454] = 8'd0;
      buffer[455] = 8'd0;
      buffer[456] = 8'd0;
      buffer[457] = 8'd0;
      buffer[458] = 8'd0;
      buffer[459] = 8'd0;
      buffer[460] = 8'd63;
      buffer[461] = 8'd128;
      buffer[462] = 8'd0;
      buffer[463] = 8'd0;
      buffer[464] = 8'd63;
      buffer[465] = 8'd128;
      buffer[466] = 8'd0;
      buffer[467] = 8'd0;
      buffer[468] = 8'd67;
      buffer[469] = 8'd122;
      buffer[470] = 8'd0;
      buffer[471] = 8'd0;
      buffer[472] = 8'd0;
      buffer[473] = 8'd0;
      buffer[474] = 8'd0;
      buffer[475] = 8'd0;
      buffer[476] = 8'd67;
      buffer[477] = 8'd83;
      buffer[478] = 8'd0;
      buffer[479] = 8'd0;
      buffer[480] = 8'd67;
      buffer[481] = 8'd83;
      buffer[482] = 8'd0;
      buffer[483] = 8'd0;
      buffer[484] = 8'd0;
      buffer[485] = 8'd0;
      buffer[486] = 8'd0;
      buffer[487] = 8'd0;
      buffer[488] = 8'd0;
      buffer[489] = 8'd0;
      buffer[490] = 8'd0;
      buffer[491] = 8'd3;
      buffer[492] = 8'd0;
      buffer[493] = 8'd0;
      buffer[494] = 8'd0;
      buffer[495] = 8'd1;
      buffer[496] = 8'd0;
      buffer[497] = 8'd0;
      buffer[498] = 8'd0;
      buffer[499] = 8'd0;
      buffer[500] = 8'd0;
      buffer[501] = 8'd0;
      buffer[502] = 8'd0;
      buffer[503] = 8'd0;
      buffer[504] = 8'd65;
      buffer[505] = 8'd112;
      buffer[506] = 8'd0;
      buffer[507] = 8'd0;
      buffer[508] = 8'd65;
      buffer[509] = 8'd112;
      buffer[510] = 8'd0;
      buffer[511] = 8'd0;
      buffer[512] = 8'd0;
      buffer[513] = 8'd0;
      buffer[514] = 8'd0;
      buffer[515] = 8'd0;
      buffer[516] = 8'd192;
      buffer[517] = 8'd160;
      buffer[518] = 8'd0;
      buffer[519] = 8'd0;
      buffer[520] = 8'd0;
      buffer[521] = 8'd0;
      buffer[522] = 8'd0;
      buffer[523] = 8'd0;
      buffer[524] = 8'd191;
      buffer[525] = 8'd128;
      buffer[526] = 8'd0;
      buffer[527] = 8'd0;
      buffer[528] = 8'd63;
      buffer[529] = 8'd128;
      buffer[530] = 8'd0;
      buffer[531] = 8'd0;
      buffer[532] = 8'd67;
      buffer[533] = 8'd122;
      buffer[534] = 8'd0;
      buffer[535] = 8'd0;
      buffer[536] = 8'd0;
      buffer[537] = 8'd0;
      buffer[538] = 8'd0;
      buffer[539] = 8'd0;
      buffer[540] = 8'd67;
      buffer[541] = 8'd83;
      buffer[542] = 8'd0;
      buffer[543] = 8'd0;
      buffer[544] = 8'd67;
      buffer[545] = 8'd83;
      buffer[546] = 8'd0;
      buffer[547] = 8'd0;
      buffer[548] = 8'd0;
      buffer[549] = 8'd0;
      buffer[550] = 8'd0;
      buffer[551] = 8'd0;
      buffer[552] = 8'd0;
      buffer[553] = 8'd0;
      buffer[554] = 8'd0;
      buffer[555] = 8'd3;
      buffer[556] = 8'd0;
      buffer[557] = 8'd0;
      buffer[558] = 8'd0;
      buffer[559] = 8'd1;
      buffer[560] = 8'd0;
      buffer[561] = 8'd0;
      buffer[562] = 8'd0;
      buffer[563] = 8'd0;
      buffer[564] = 8'd65;
      buffer[565] = 8'd112;
      buffer[566] = 8'd0;
      buffer[567] = 8'd0;
      buffer[568] = 8'd65;
      buffer[569] = 8'd200;
      buffer[570] = 8'd0;
      buffer[571] = 8'd0;
      buffer[572] = 8'd65;
      buffer[573] = 8'd200;
      buffer[574] = 8'd0;
      buffer[575] = 8'd0;
      buffer[576] = 8'd0;
      buffer[577] = 8'd0;
      buffer[578] = 8'd0;
      buffer[579] = 8'd0;
      buffer[580] = 8'd192;
      buffer[581] = 8'd160;
      buffer[582] = 8'd0;
      buffer[583] = 8'd0;
      buffer[584] = 8'd66;
      buffer[585] = 8'd140;
      buffer[586] = 8'd0;
      buffer[587] = 8'd0;
      buffer[588] = 8'd63;
      buffer[589] = 8'd128;
      buffer[590] = 8'd0;
      buffer[591] = 8'd0;
      buffer[592] = 8'd63;
      buffer[593] = 8'd128;
      buffer[594] = 8'd0;
      buffer[595] = 8'd0;
      buffer[596] = 8'd67;
      buffer[597] = 8'd122;
      buffer[598] = 8'd0;
      buffer[599] = 8'd0;
      buffer[600] = 8'd67;
      buffer[601] = 8'd83;
      buffer[602] = 8'd0;
      buffer[603] = 8'd0;
      buffer[604] = 8'd0;
      buffer[605] = 8'd0;
      buffer[606] = 8'd0;
      buffer[607] = 8'd0;
      buffer[608] = 8'd0;
      buffer[609] = 8'd0;
      buffer[610] = 8'd0;
      buffer[611] = 8'd0;
      buffer[612] = 8'd0;
      buffer[613] = 8'd0;
      buffer[614] = 8'd0;
      buffer[615] = 8'd0;
      buffer[616] = 8'd0;
      buffer[617] = 8'd0;
      buffer[618] = 8'd0;
      buffer[619] = 8'd1;
      buffer[620] = 8'd0;
      buffer[621] = 8'd0;
      buffer[622] = 8'd0;
      buffer[623] = 8'd1;
      buffer[624] = 8'd0;
      buffer[625] = 8'd0;
      buffer[626] = 8'd0;
      buffer[627] = 8'd0;
      buffer[628] = 8'd64;
      buffer[629] = 8'd160;
      buffer[630] = 8'd0;
      buffer[631] = 8'd0;
      buffer[632] = 8'd65;
      buffer[633] = 8'd48;
      buffer[634] = 8'd0;
      buffer[635] = 8'd0;
      buffer[636] = 8'd66;
      buffer[637] = 8'd52;
      buffer[638] = 8'd0;
      buffer[639] = 8'd0;
      buffer[640] = 8'd0;
      buffer[641] = 8'd0;
      buffer[642] = 8'd0;
      buffer[643] = 8'd0;
      buffer[644] = 8'd66;
      buffer[645] = 8'd12;
      buffer[646] = 8'd0;
      buffer[647] = 8'd0;
      buffer[648] = 8'd66;
      buffer[649] = 8'd32;
      buffer[650] = 8'd0;
      buffer[651] = 8'd0;
      buffer[652] = 8'd63;
      buffer[653] = 8'd128;
      buffer[654] = 8'd0;
      buffer[655] = 8'd0;
      buffer[656] = 8'd63;
      buffer[657] = 8'd128;
      buffer[658] = 8'd0;
      buffer[659] = 8'd0;
      buffer[660] = 8'd67;
      buffer[661] = 8'd122;
      buffer[662] = 8'd0;
      buffer[663] = 8'd0;
      buffer[664] = 8'd67;
      buffer[665] = 8'd83;
      buffer[666] = 8'd0;
      buffer[667] = 8'd0;
      buffer[668] = 8'd67;
      buffer[669] = 8'd0;
      buffer[670] = 8'd0;
      buffer[671] = 8'd0;
      buffer[672] = 8'd0;
      buffer[673] = 8'd0;
      buffer[674] = 8'd0;
      buffer[675] = 8'd0;
      buffer[676] = 8'd0;
      buffer[677] = 8'd0;
      buffer[678] = 8'd0;
      buffer[679] = 8'd0;
      buffer[680] = 8'd0;
      buffer[681] = 8'd0;
      buffer[682] = 8'd0;
      buffer[683] = 8'd3;
      buffer[684] = 8'd0;
      buffer[685] = 8'd0;
      buffer[686] = 8'd0;
      buffer[687] = 8'd1;
      buffer[688] = 8'd0;
      buffer[689] = 8'd0;
      buffer[690] = 8'd0;
      buffer[691] = 8'd0;
      buffer[692] = 8'd65;
      buffer[693] = 8'd240;
      buffer[694] = 8'd0;
      buffer[695] = 8'd0;
      buffer[696] = 8'd66;
      buffer[697] = 8'd52;
      buffer[698] = 8'd0;
      buffer[699] = 8'd0;
      buffer[700] = 8'd66;
      buffer[701] = 8'd150;
      buffer[702] = 8'd0;
      buffer[703] = 8'd0;
      buffer[704] = 8'd0;
      buffer[705] = 8'd0;
      buffer[706] = 8'd0;
      buffer[707] = 8'd0;
      buffer[708] = 8'd0;
      buffer[709] = 8'd0;
      buffer[710] = 8'd0;
      buffer[711] = 8'd0;
      buffer[712] = 8'd66;
      buffer[713] = 8'd32;
      buffer[714] = 8'd0;
      buffer[715] = 8'd0;
      buffer[716] = 8'd63;
      buffer[717] = 8'd128;
      buffer[718] = 8'd0;
      buffer[719] = 8'd0;
      buffer[720] = 8'd63;
      buffer[721] = 8'd128;
      buffer[722] = 8'd0;
      buffer[723] = 8'd0;
      buffer[724] = 8'd67;
      buffer[725] = 8'd122;
      buffer[726] = 8'd0;
      buffer[727] = 8'd0;
      buffer[728] = 8'd67;
      buffer[729] = 8'd83;
      buffer[730] = 8'd0;
      buffer[731] = 8'd0;
      buffer[732] = 8'd67;
      buffer[733] = 8'd0;
      buffer[734] = 8'd0;
      buffer[735] = 8'd0;
      buffer[736] = 8'd0;
      buffer[737] = 8'd0;
      buffer[738] = 8'd0;
      buffer[739] = 8'd0;
      buffer[740] = 8'd0;
      buffer[741] = 8'd0;
      buffer[742] = 8'd0;
      buffer[743] = 8'd0;
      buffer[744] = 8'd0;
      buffer[745] = 8'd0;
      buffer[746] = 8'd0;
      buffer[747] = 8'd1;
      buffer[748] = 8'd0;
      buffer[749] = 8'd0;
      buffer[750] = 8'd0;
      buffer[751] = 8'd1;
      buffer[752] = 8'd0;
      buffer[753] = 8'd0;
      buffer[754] = 8'd0;
      buffer[755] = 8'd0;
      buffer[756] = 8'd65;
      buffer[757] = 8'd200;
      buffer[758] = 8'd0;
      buffer[759] = 8'd0;
      buffer[760] = 8'd66;
      buffer[761] = 8'd36;
      buffer[762] = 8'd0;
      buffer[763] = 8'd0;
      buffer[764] = 8'd66;
      buffer[765] = 8'd140;
      buffer[766] = 8'd0;
      buffer[767] = 8'd0;
      buffer[768] = 8'd0;
      buffer[769] = 8'd0;
      buffer[770] = 8'd0;
      buffer[771] = 8'd0;
      buffer[772] = 8'd64;
      buffer[773] = 8'd160;
      buffer[774] = 8'd0;
      buffer[775] = 8'd0;
      buffer[776] = 8'd66;
      buffer[777] = 8'd32;
      buffer[778] = 8'd0;
      buffer[779] = 8'd0;
      buffer[780] = 8'd63;
      buffer[781] = 8'd128;
      buffer[782] = 8'd0;
      buffer[783] = 8'd0;
      buffer[784] = 8'd63;
      buffer[785] = 8'd128;
      buffer[786] = 8'd0;
      buffer[787] = 8'd0;
      buffer[788] = 8'd67;
      buffer[789] = 8'd122;
      buffer[790] = 8'd0;
      buffer[791] = 8'd0;
      buffer[792] = 8'd0;
      buffer[793] = 8'd0;
      buffer[794] = 8'd0;
      buffer[795] = 8'd0;
      buffer[796] = 8'd0;
      buffer[797] = 8'd0;
      buffer[798] = 8'd0;
      buffer[799] = 8'd0;
      buffer[800] = 8'd0;
      buffer[801] = 8'd0;
      buffer[802] = 8'd0;
      buffer[803] = 8'd0;
      buffer[804] = 8'd0;
      buffer[805] = 8'd0;
      buffer[806] = 8'd0;
      buffer[807] = 8'd1;
      buffer[808] = 8'd0;
      buffer[809] = 8'd0;
      buffer[810] = 8'd0;
      buffer[811] = 8'd1;
      buffer[812] = 8'd0;
      buffer[813] = 8'd0;
      buffer[814] = 8'd0;
      buffer[815] = 8'd1;
      buffer[816] = 8'd0;
      buffer[817] = 8'd0;
      buffer[818] = 8'd0;
      buffer[819] = 8'd0;
      buffer[820] = 8'd66;
      buffer[821] = 8'd200;
      buffer[822] = 8'd0;
      buffer[823] = 8'd0;
      buffer[824] = 8'd64;
      buffer[825] = 8'd160;
      buffer[826] = 8'd0;
      buffer[827] = 8'd0;
      buffer[828] = 8'd67;
      buffer[829] = 8'd72;
      buffer[830] = 8'd0;
      buffer[831] = 8'd0;
      buffer[832] = 8'd0;
      buffer[833] = 8'd0;
      buffer[834] = 8'd0;
      buffer[835] = 8'd0;
      buffer[836] = 8'd194;
      buffer[837] = 8'd12;
      buffer[838] = 8'd0;
      buffer[839] = 8'd0;
      buffer[840] = 8'd67;
      buffer[841] = 8'd22;
      buffer[842] = 8'd0;
      buffer[843] = 8'd0;
      buffer[844] = 8'd63;
      buffer[845] = 8'd128;
      buffer[846] = 8'd0;
      buffer[847] = 8'd0;
      buffer[848] = 8'd63;
      buffer[849] = 8'd128;
      buffer[850] = 8'd0;
      buffer[851] = 8'd0;
      buffer[852] = 8'd67;
      buffer[853] = 8'd122;
      buffer[854] = 8'd0;
      buffer[855] = 8'd0;
      buffer[856] = 8'd67;
      buffer[857] = 8'd72;
      buffer[858] = 8'd0;
      buffer[859] = 8'd0;
      buffer[860] = 8'd67;
      buffer[861] = 8'd72;
      buffer[862] = 8'd0;
      buffer[863] = 8'd0;
      buffer[864] = 8'd67;
      buffer[865] = 8'd72;
      buffer[866] = 8'd0;
      buffer[867] = 8'd0;
      buffer[868] = 8'd0;
      buffer[869] = 8'd0;
      buffer[870] = 8'd0;
      buffer[871] = 8'd0;
      buffer[872] = 8'd0;
      buffer[873] = 8'd0;
      buffer[874] = 8'd0;
      buffer[875] = 8'd3;
      buffer[876] = 8'd0;
      buffer[877] = 8'd0;
      buffer[878] = 8'd0;
      buffer[879] = 8'd1;
      buffer[880] = 8'd0;
      buffer[881] = 8'd0;
      buffer[882] = 8'd0;
      buffer[883] = 8'd0;
      buffer[884] = 8'd65;
      buffer[885] = 8'd200;
      buffer[886] = 8'd0;
      buffer[887] = 8'd0;
      buffer[888] = 8'd65;
      buffer[889] = 8'd32;
      buffer[890] = 8'd0;
      buffer[891] = 8'd0;
      buffer[892] = 8'd65;
      buffer[893] = 8'd32;
      buffer[894] = 8'd0;
      buffer[895] = 8'd0;
      buffer[896] = 8'd0;
      buffer[897] = 8'd0;
      buffer[898] = 8'd0;
      buffer[899] = 8'd0;
      buffer[900] = 8'd192;
      buffer[901] = 8'd160;
      buffer[902] = 8'd0;
      buffer[903] = 8'd0;
      buffer[904] = 8'd0;
      buffer[905] = 8'd0;
      buffer[906] = 8'd0;
      buffer[907] = 8'd0;
      buffer[908] = 8'd63;
      buffer[909] = 8'd128;
      buffer[910] = 8'd0;
      buffer[911] = 8'd0;
      buffer[912] = 8'd63;
      buffer[913] = 8'd128;
      buffer[914] = 8'd0;
      buffer[915] = 8'd0;
      buffer[916] = 8'd67;
      buffer[917] = 8'd122;
      buffer[918] = 8'd0;
      buffer[919] = 8'd0;
      buffer[920] = 8'd67;
      buffer[921] = 8'd83;
      buffer[922] = 8'd0;
      buffer[923] = 8'd0;
      buffer[924] = 8'd67;
      buffer[925] = 8'd0;
      buffer[926] = 8'd0;
      buffer[927] = 8'd0;
      buffer[928] = 8'd67;
      buffer[929] = 8'd0;
      buffer[930] = 8'd0;
      buffer[931] = 8'd0;
      buffer[932] = 8'd0;
      buffer[933] = 8'd0;
      buffer[934] = 8'd0;
      buffer[935] = 8'd0;
      buffer[936] = 8'd0;
      buffer[937] = 8'd0;
      buffer[938] = 8'd0;
      buffer[939] = 8'd3;
      buffer[940] = 8'd0;
      buffer[941] = 8'd0;
      buffer[942] = 8'd0;
      buffer[943] = 8'd2;
      buffer[944] = 8'd0;
      buffer[945] = 8'd0;
      buffer[946] = 8'd0;
      buffer[947] = 8'd0;
      buffer[948] = 8'd65;
      buffer[949] = 8'd200;
      buffer[950] = 8'd0;
      buffer[951] = 8'd0;
      buffer[952] = 8'd65;
      buffer[953] = 8'd160;
      buffer[954] = 8'd0;
      buffer[955] = 8'd0;
      buffer[956] = 8'd65;
      buffer[957] = 8'd160;
      buffer[958] = 8'd0;
      buffer[959] = 8'd0;
      buffer[960] = 8'd0;
      buffer[961] = 8'd0;
      buffer[962] = 8'd0;
      buffer[963] = 8'd0;
      buffer[964] = 8'd0;
      buffer[965] = 8'd0;
      buffer[966] = 8'd0;
      buffer[967] = 8'd0;
      buffer[968] = 8'd66;
      buffer[969] = 8'd140;
      buffer[970] = 8'd0;
      buffer[971] = 8'd0;
      buffer[972] = 8'd63;
      buffer[973] = 8'd128;
      buffer[974] = 8'd0;
      buffer[975] = 8'd0;
      buffer[976] = 8'd62;
      buffer[977] = 8'd153;
      buffer[978] = 8'd153;
      buffer[979] = 8'd154;
      buffer[980] = 8'd0;
      buffer[981] = 8'd0;
      buffer[982] = 8'd0;
      buffer[983] = 8'd0;
      buffer[984] = 8'd0;
      buffer[985] = 8'd0;
      buffer[986] = 8'd0;
      buffer[987] = 8'd0;
      buffer[988] = 8'd0;
      buffer[989] = 8'd0;
      buffer[990] = 8'd0;
      buffer[991] = 8'd0;
      buffer[992] = 8'd67;
      buffer[993] = 8'd127;
      buffer[994] = 8'd0;
      buffer[995] = 8'd0;
      buffer[996] = 8'd0;
      buffer[997] = 8'd0;
      buffer[998] = 8'd0;
      buffer[999] = 8'd2;
      buffer[1000] = 8'd0;
      buffer[1001] = 8'd0;
      buffer[1002] = 8'd0;
      buffer[1003] = 8'd3;
      buffer[1004] = 8'd0;
      buffer[1005] = 8'd0;
      buffer[1006] = 8'd0;
      buffer[1007] = 8'd1;
      buffer[1008] = 8'd0;
      buffer[1009] = 8'd0;
      buffer[1010] = 8'd0;
      buffer[1011] = 8'd0;
      buffer[1012] = 8'd65;
      buffer[1013] = 8'd160;
      buffer[1014] = 8'd0;
      buffer[1015] = 8'd0;
      buffer[1016] = 8'd65;
      buffer[1017] = 8'd160;
      buffer[1018] = 8'd0;
      buffer[1019] = 8'd0;
      buffer[1020] = 8'd65;
      buffer[1021] = 8'd160;
      buffer[1022] = 8'd0;
      buffer[1023] = 8'd0;
      buffer[1024] = 8'd66;
      buffer[1025] = 8'd200;
      buffer[1026] = 8'd0;
      buffer[1027] = 8'd0;
      buffer[1028] = 8'd66;
      buffer[1029] = 8'd32;
      buffer[1030] = 8'd0;
      buffer[1031] = 8'd0;
      buffer[1032] = 8'd66;
      buffer[1033] = 8'd240;
      buffer[1034] = 8'd0;
      buffer[1035] = 8'd0;
      buffer[1036] = 8'd63;
      buffer[1037] = 8'd128;
      buffer[1038] = 8'd0;
      buffer[1039] = 8'd0;
      buffer[1040] = 8'd63;
      buffer[1041] = 8'd128;
      buffer[1042] = 8'd0;
      buffer[1043] = 8'd0;
      buffer[1044] = 8'd67;
      buffer[1045] = 8'd22;
      buffer[1046] = 8'd0;
      buffer[1047] = 8'd0;
      buffer[1048] = 8'd67;
      buffer[1049] = 8'd127;
      buffer[1050] = 8'd0;
      buffer[1051] = 8'd0;
      buffer[1052] = 8'd67;
      buffer[1053] = 8'd127;
      buffer[1054] = 8'd0;
      buffer[1055] = 8'd0;
      buffer[1056] = 8'd67;
      buffer[1057] = 8'd127;
      buffer[1058] = 8'd0;
      buffer[1059] = 8'd0;
      buffer[1060] = 8'd0;
      buffer[1061] = 8'd0;
      buffer[1062] = 8'd0;
      buffer[1063] = 8'd0;
      buffer[1064] = 8'd0;
      buffer[1065] = 8'd0;
      buffer[1066] = 8'd0;
      buffer[1067] = 8'd2;
      buffer[1068] = 8'd0;
      buffer[1069] = 8'd0;
      buffer[1070] = 8'd0;
      buffer[1071] = 8'd2;
      buffer[1072] = 8'd0;
      buffer[1073] = 8'd0;
      buffer[1074] = 8'd0;
      buffer[1075] = 8'd0;
      buffer[1076] = 8'd0;
      buffer[1077] = 8'd0;
      buffer[1078] = 8'd0;
      buffer[1079] = 8'd0;
      buffer[1080] = 8'd0;
      buffer[1081] = 8'd0;
      buffer[1082] = 8'd0;
      buffer[1083] = 8'd0;
      buffer[1084] = 8'd191;
      buffer[1085] = 8'd128;
      buffer[1086] = 8'd0;
      buffer[1087] = 8'd0;
      buffer[1088] = 8'd0;
      buffer[1089] = 8'd0;
      buffer[1090] = 8'd0;
      buffer[1091] = 8'd0;
      buffer[1092] = 8'd0;
      buffer[1093] = 8'd0;
      buffer[1094] = 8'd0;
      buffer[1095] = 8'd0;
      buffer[1096] = 8'd67;
      buffer[1097] = 8'd72;
      buffer[1098] = 8'd0;
      buffer[1099] = 8'd0;
      buffer[1100] = 8'd63;
      buffer[1101] = 8'd128;
      buffer[1102] = 8'd0;
      buffer[1103] = 8'd0;
      buffer[1104] = 8'd62;
      buffer[1105] = 8'd76;
      buffer[1106] = 8'd204;
      buffer[1107] = 8'd205;
      buffer[1108] = 8'd0;
      buffer[1109] = 8'd0;
      buffer[1110] = 8'd0;
      buffer[1111] = 8'd0;
      buffer[1112] = 8'd67;
      buffer[1113] = 8'd127;
      buffer[1114] = 8'd0;
      buffer[1115] = 8'd0;
      buffer[1116] = 8'd0;
      buffer[1117] = 8'd0;
      buffer[1118] = 8'd0;
      buffer[1119] = 8'd0;
      buffer[1120] = 8'd0;
      buffer[1121] = 8'd0;
      buffer[1122] = 8'd0;
      buffer[1123] = 8'd0;
      buffer[1124] = 8'd255;
      buffer[1125] = 8'd255;
      buffer[1126] = 8'd255;
      buffer[1127] = 8'd255;
      buffer[1128] = 8'd0;
      buffer[1129] = 8'd0;
      buffer[1130] = 8'd0;
      buffer[1131] = 8'd0;
      buffer[1132] = 8'd0;
      buffer[1133] = 8'd0;
      buffer[1134] = 8'd0;
      buffer[1135] = 8'd1;
      buffer[1136] = 8'd0;
      buffer[1137] = 8'd0;
      buffer[1138] = 8'd0;
      buffer[1139] = 8'd2;
      buffer[1140] = 8'd255;
      buffer[1141] = 8'd255;
      buffer[1142] = 8'd255;
      buffer[1143] = 8'd255;
      buffer[1144] = 8'd0;
      buffer[1145] = 8'd0;
      buffer[1146] = 8'd0;
      buffer[1147] = 8'd3;
      buffer[1148] = 8'd0;
      buffer[1149] = 8'd0;
      buffer[1150] = 8'd0;
      buffer[1151] = 8'd1;
      buffer[1152] = 8'd0;
      buffer[1153] = 8'd0;
      buffer[1154] = 8'd0;
      buffer[1155] = 8'd4;
      buffer[1156] = 8'd255;
      buffer[1157] = 8'd255;
      buffer[1158] = 8'd255;
      buffer[1159] = 8'd255;
      buffer[1160] = 8'd0;
      buffer[1161] = 8'd0;
      buffer[1162] = 8'd0;
      buffer[1163] = 8'd5;
      buffer[1164] = 8'd0;
      buffer[1165] = 8'd0;
      buffer[1166] = 8'd0;
      buffer[1167] = 8'd6;
      buffer[1168] = 8'd0;
      buffer[1169] = 8'd0;
      buffer[1170] = 8'd0;
      buffer[1171] = 8'd7;
      buffer[1172] = 8'd255;
      buffer[1173] = 8'd255;
      buffer[1174] = 8'd255;
      buffer[1175] = 8'd255;
      buffer[1176] = 8'd0;
      buffer[1177] = 8'd0;
      buffer[1178] = 8'd0;
      buffer[1179] = 8'd8;
      buffer[1180] = 8'd255;
      buffer[1181] = 8'd255;
      buffer[1182] = 8'd255;
      buffer[1183] = 8'd255;
      buffer[1184] = 8'd0;
      buffer[1185] = 8'd0;
      buffer[1186] = 8'd0;
      buffer[1187] = 8'd9;
      buffer[1188] = 8'd0;
      buffer[1189] = 8'd0;
      buffer[1190] = 8'd0;
      buffer[1191] = 8'd10;
      buffer[1192] = 8'd255;
      buffer[1193] = 8'd255;
      buffer[1194] = 8'd255;
      buffer[1195] = 8'd255;
      buffer[1196] = 8'd0;
      buffer[1197] = 8'd0;
      buffer[1198] = 8'd0;
      buffer[1199] = 8'd12;
      buffer[1200] = 8'd255;
      buffer[1201] = 8'd255;
      buffer[1202] = 8'd255;
      buffer[1203] = 8'd255;
      buffer[1204] = 8'd0;
      buffer[1205] = 8'd0;
      buffer[1206] = 8'd0;
      buffer[1207] = 8'd13;
      buffer[1208] = 8'd255;
      buffer[1209] = 8'd255;
      buffer[1210] = 8'd255;
      buffer[1211] = 8'd255;
      buffer[1212] = 8'd0;
      buffer[1213] = 8'd0;
      buffer[1214] = 8'd0;
      buffer[1215] = 8'd14;
      buffer[1216] = 8'd255;
      buffer[1217] = 8'd255;
      buffer[1218] = 8'd255;
      buffer[1219] = 8'd255;
      buffer[1220] = 8'd0;
      buffer[1221] = 8'd0;
      buffer[1222] = 8'd0;
      buffer[1223] = 8'd15;
      buffer[1224] = 8'd255;
      buffer[1225] = 8'd255;
      buffer[1226] = 8'd255;
      buffer[1227] = 8'd255;
      buffer[1228] = 8'd0;
      buffer[1229] = 8'd0;
      buffer[1230] = 8'd0;
      buffer[1231] = 8'd16;
      buffer[1232] = 8'd255;
      buffer[1233] = 8'd255;
      buffer[1234] = 8'd255;
      buffer[1235] = 8'd255;
      buffer[1236] = 8'd255;
      buffer[1237] = 8'd255;
      buffer[1238] = 8'd255;
      buffer[1239] = 8'd255;
      buffer[1240] = 8'd0;
      buffer[1241] = 8'd0;
      buffer[1242] = 8'd0;
      buffer[1243] = 8'd11;
      buffer[1244] = 8'd0;
      buffer[1245] = 8'd0;
      buffer[1246] = 8'd0;
      buffer[1247] = 8'd0;
      buffer[1248] = 8'd0;
      buffer[1249] = 8'd0;
      buffer[1250] = 8'd0;
      buffer[1251] = 8'd1;
      buffer[1252] = 8'd0;
      buffer[1253] = 8'd0;
      buffer[1254] = 8'd0;
      buffer[1255] = 8'd2;
      buffer[1256] = 8'd0;
      buffer[1257] = 8'd0;
      buffer[1258] = 8'd0;
      buffer[1259] = 8'd3;
      buffer[1260] = 8'd0;
      buffer[1261] = 8'd0;
      buffer[1262] = 8'd0;
      buffer[1263] = 8'd4;
      buffer[1264] = 8'd0;
      buffer[1265] = 8'd0;
      buffer[1266] = 8'd0;
      buffer[1267] = 8'd6;
      buffer[1268] = 8'd255;
      buffer[1269] = 8'd255;
      buffer[1270] = 8'd255;
      buffer[1271] = 8'd255;
      buffer[1272] = 8'd0;
      buffer[1273] = 8'd0;
      buffer[1274] = 8'd0;
      buffer[1275] = 8'd99;
      buffer[1276] = 8'd0;
      buffer[1277] = 8'd0;
      buffer[1278] = 8'd0;
      buffer[1279] = 8'd9;
      buffer[1280] = 8'd0;
      buffer[1281] = 8'd0;
      buffer[1282] = 8'd0;
      buffer[1283] = 8'd8;
      buffer[1284] = 8'd0;
      buffer[1285] = 8'd0;
      buffer[1286] = 8'd0;
      buffer[1287] = 8'd7;
      buffer[1288] = 8'd0;
      buffer[1289] = 8'd0;
      buffer[1290] = 8'd0;
      buffer[1291] = 8'd5;
      buffer[1292] = 8'd255;
      buffer[1293] = 8'd255;
      buffer[1294] = 8'd255;
      buffer[1295] = 8'd255;
      buffer[1296] = 8'd255;
      buffer[1297] = 8'd255;
      buffer[1298] = 8'd255;
      buffer[1299] = 8'd255;
   end // initial begin

   
   // Reply to MMU
   /////////////
   reg [3:0] addr_cache;      
   always @(posedge clk) begin
      if(rstn) begin
         if (reading_state == r_waiting_ready) begin
            if (mmu_axi_arvalid) begin
               mmu_axi_arready <= 0;               
               if(mmu_axi_araddr[3:0] == 4'h0 && !is_buffer_empty) begin
                  mmu_axi_rvalid <= 1;
                  head_idx <= head_idx + 1;                  
                  mmu_axi_rdata <= {24'b0, buffer[head_idx]};
                  mmu_axi_rresp <= 2'b00;                  
                  reading_state <= r_writing_data;                  
               end else begin                              
                  uart_axi_arvalid <= 1;
                  uart_axi_araddr <= mmu_axi_araddr[3:0];
                  addr_cache <= mmu_axi_araddr[3:0];
                  uart_axi_arprot <= mmu_axi_arprot;                                    
                  reading_state <= r_writing_ready;
               end               
            end else begin
               mmu_axi_arready <= 0;
               uart_axi_arvalid <= 1;
               uart_axi_araddr <= 4'b0;
               uart_axi_arprot <= 3'b0;               
               reading_state <= r_waiting_uartlite_arready;
            end
         end else if (reading_state == r_writing_ready) begin
            if(uart_axi_arready) begin
               uart_axi_arvalid <= 0;            
               uart_axi_rready <= 1;            
               reading_state <= r_waiting_data;
            end
         end if (reading_state == r_waiting_data) begin
            if (uart_axi_rvalid) begin
               uart_axi_rready <= 0;
               mmu_axi_rvalid <= 1;
               if (addr_cache == 4'h8) begin
                  mmu_axi_rdata <= {uart_axi_rdata[31:1], !is_buffer_empty | uart_axi_rdata[0]};
               end else begin
                  mmu_axi_rdata <= uart_axi_rdata;
               end
               mmu_axi_rresp <= uart_axi_rresp;   
               reading_state <= r_writing_data;            
            end
         end if (reading_state == r_writing_data) begin
            if(mmu_axi_rready) begin
               mmu_axi_rvalid <= 0;
               mmu_axi_arready <= 1;
               reading_state <= r_waiting_ready;
            end
         end if (reading_state == r_waiting_uartlite_arready) begin
            if(uart_axi_arready) begin
               uart_axi_arvalid <= 0;            
               uart_axi_rready <= 1;            
               reading_state <= r_waiting_uartlite_rvalid;               
            end
         end if (reading_state == r_waiting_uartlite_rvalid) begin
            if (uart_axi_rvalid) begin
               uart_axi_rready <= 0;
               if (uart_axi_rresp == 2'b00) begin
                  // if valid data exists
                  buffer[tail_idx] <= uart_axi_rdata[7:0];
                  tail_idx <= tail_idx + 1;
               end
               mmu_axi_arready <= 1;
               reading_state <= r_waiting_ready;            
            end
         end
      end
   end      
endmodule
`default_nettype wire
