typedef struct packed {
   logic addi;   
   logic add;
   logic beq;
   logic jal;
} instructions;
